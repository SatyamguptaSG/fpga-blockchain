module com8bit(a[7:0],b[7:0],alb,aeb,agb);
assign agb=(a[7]&(a[7]^b[7]))^(a[6]&(a[6]^b[6]))^(a[5]&(a[5]^b[5]))^(a[4]&(a[4]^b[4]))^(a[3]&(a[3]^b[3]))^(a[2]&(a[2]^b[2]))^(a[1]&(a[1]^b[1]))^(a[0]&(a[0]^b[0]))
assign alb=(b[7]&(a[7]^b[7]))^(b[6]&(a[6]^b[6]))^(b[5]&(a[5]^b[5]))^(b[4]&(a[4]^b[4]))^(b[3]&(a[3]^b[3]))^(b[2]&(a[2]^b[2]))^(b[1]&(a[1]^b[1]))^(b[0]&(a[0]^b[0]))
assign aeb=(a[7]&b[7])&(a[6]&b[6])&(a[5]&b[5])&(a[4]&b[4])&(a[3]&b[3])&(a[2]&b[2])&(a[1]&b[1])&(a[0]&b[0])
endmodule
